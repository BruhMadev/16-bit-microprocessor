`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.09.2021 08:55:21
// Design Name: 
// Module Name: alu_control_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_control_unit(
// takes parts of the instruction (funct) and part of controll signal generated by control_unit (alu_op) 
// and generates corresponding signal for ALU to ADD, SUB,, AND, OR or compare. 
input [1:0] alu_op, input [3:0] funct, output reg [2:0] ALU_control, output JR_control
    );
    wire [5:0]ALU_control_in;
    assign ALU_control_in = {alu_op, funct};
    always@(ALU_control_in)
    begin
    casex (ALU_control_in)
    6'b11xxxx: ALU_control = 3'b000; // add (for addi LW and SW) I-type
    6'b10xxxx: ALU_control = 3'b100; // compare (for slti) I-type
    6'b01xxxx: ALU_control = 3'b001; // sub (for beq) if they are equal alu outputs 0, I-type
    6'b000000: ALU_control = 3'b000; // add for, R-type add funct = 4'b0 
    6'b000001: ALU_control = 3'b001; // sub for Rtype 
    6'b000010: ALU_control = 3'b010; // and   
    6'b000011: ALU_control = 3'b011; // OR
    6'b000100: ALU_control = 3'b100; // compare (strictly less than)
    default: ALU_control = 3'b000;
    endcase
    end
    assign JR_control = (ALU_control_in == 6'b001000) ? 1'b1 : 1'b0;
endmodule
